B
0 0 0 0 0 r h 1 B 8 B
0 0 0 0 0 r h 2 B 7 B
0 0 0 0 0 r h 3 B 6 B
0 0 0 0 0 r h 4 B 5 B
4 11 1 2 2 12 1 10 1 4 3 5 4 8 5 7 0 10 1 4 3 11 4 9 0 5 0 6 2 6 2 3 3 3 0 9 2 8
